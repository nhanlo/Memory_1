`define lb  3'h000
`define lh  3'h010
`define lbu 3'h100
`define lhu 3'h110
`define sb  3'h001

